 

`uvm_info("FINAL_PHASE_TOPDOWN"," FINAL_PHASE   IS STARTED ",UVM_NONE)

`uvm_info("FINAL_PHASE_TOPDOWN"," FINAL_PHASE  IS ENDED ",UVM_NONE)